BZh91AY&SY~���߀ryg����߰?���a� ����	l��P�\��T��k�,�-��SF���PUSY � ��@��6kZ�m���    �>��#QJ;�9�Õ�(J���3��w�z�ڥJ�����T����y"���ֹ@*��V�*��@Q@ ���-� R�||�
(QW��EO��9��+Z4�ܡ2i(S�E��(W��>��[�P��mc���\cl�e���������+M�F�7��X�tu��T)JX�(�Q��l�Z�ݕ�����2ik�\6X����=�J����l�3>#�lf�67N��ۍhmeZgg8�ڊ���ȥJ�UJc���k�6jl3c�y��8��6L�gv�=�Tw����B!}@�QQ��{��ǜ�cB���W��NW.�k5�=����B�[�J@Q_}�ۏmX|��m����w���� �kU��غr��&�Z�h���'�!��)��-��y�M��5���OYҍ�-�1��t�W��Ͼ���AI�z��Y|�[Y���摃)Ev����=ή��v$�m2h E���,<Q{쭾�m�xx8�l�+[����Qn��Y���@  �(� � *�       	T��J�M0�d�� 0!���DR*(�00 C �ɀ%M����OD`�L�M#!�4 d� Jz&����ѓ&F��2b4��bi��L�iH1�&�٩6Ҟ��O	JR�@0�@��� �4��>���$��	3�  )����p���� �'���0���j���E@R����O����~�)��N�TTM�
8?��sܞ���&��ԛ���@O���?�=>�'���c>��A�Lz����`O���������X��ق��M�~���u��}��Z4��p��@S悇ȑ5�(�����OH��߹$�I$�A���ߧJ**'X� ��
 81`-"��t�OgI�BOI�R�Y�ZA]BȠ
�fz�����\�����~#���P�������b����=Hc��c���M��P ��PDU�"��@B@P?_��� �����}���]c���a���Oz|?�G���U`���_'͊���O�����`��Iͷ
7Ðz�M�nF���b��|Ƴ�B�ޠJ�1�eߨ^�	I;zm�|!�����9���ñ˱Ͳ��$)��њ���X�b#kS�b��'z�^��T{²(c��̺���M�vse0�֍��tCעqE��/�̧���b�����^F��7��F���W���EU�������z-�a�˶����3~�rlɷǅ�%���h��i�ݦp�4k��ޙS�)���5�:h�!��N7�[n(���N�����Kz��QEoMYk���X�L|�Qj&�!��8���1JU�j���Z3��ɻG��gg�5'V��E�8�U��º��ar}��`߸F{뾧�-�UE�Fr�Ί�Uy0���y����[����溮x]C�O^2��\5��{��Cc�������O�'��Uo�5V�*������G��s�nx!�a�;���}fզ��3QE'�6׍��Y�2uӄp+��%f�ܜ51�^�r�L\�&j�i��)�ǳ��2K�Ӆ��-\�ٳ��f��j|�T����g9�1D��Jf���Wx�8�T�����7CzN����a'+,oq���kfC�Qp��;�tv�k;��r-����f]��m_º��-LB�����r}z{7s�[�,��S9�Pv��ӹ�h���秝f�>��[���!;/)a}���h�NSP�qZ0��7b�q�N9f��v�t���ݬ�C�9aK��>�zO�7�[4C���n/dѸr��[�.P�a͓�p}�"��ڢ�<^��]{�P4\.�iQ�:���{9�Hl�V2�kPwXhu�|�R��}���'��S�k9|�Ff�t�ިl���9v<�+�	vWm7#0���=�墳(ly{��û�e��v�u�Y��Ŷ�O	G�D+0�3!&p��2�)��h�Q�VR��4�bN�X�,�%�b�^�����k�gH��-Z�@[o'x,��}����.�DQ�Ҙ:��5��zcY�h|���f�K.�#���)�
w���SW129��և�WWu��^��,�̴٣T���3Ν�.�42b�����7�C��N1�,F,�WM��Ɋ��j��2n^5�ʹ6ju�.�]9����͜�#���=�6G�Z-�H�y���&�ZY��O\�65�;6�~�]y���r�(`����	�����7�lGy����f���p���s�����%qF��W�vz�V�V3�b7��5���5�P�m�)�ZHg2��
��|a�E��������FP>�vR�pԼ�TY��
��.����OR��C�\�4Y�L{�T��k�0�|I�F���f�u�x������
���g�/x�r��:�f�f�Y�V|`�Qg@�{�t��MUz�3�{15���5�9�]F;�V�\Lժ�j'�]]:��f�����M��M��ިNVR�e-=,]�vY��γ�=��2h����_1Uv`л�D�(�E��YT�S{�LMi��[�
݁u�a���w͡U�%���:�A=no*��!C�-֘?#:�j�ȳ���E��c���VC�f�&YTxE��-�X�������e�]�έ�(Q�?g�2m�pѯ9��sd7iKsFcע�����a)�G�o���<yQO#�6��djSwV,��B��
C8S��⩳i�҆�Jfm�~d�Ù]��&yS&ʮ�^>U�tí�$j,�q��t��(>�o}(�8��p�̽�gi���M�v�ZZ���Oo������).�j�k��SV�a�W]�>���S���)i����3(����іm�#�Í�3y|��}�o/&4k��y=�)���5�TΒ��sE)����UG<aw�Q�
(��(��;�U��&^�/����l��u�wxE�k�K��9��ş_���DOjE��\gb]UMb�2y4h�iy_:m<#���[�F���:_I���W��f�a{�#�1�4a��x^��g���5a�a�f�a�mXџL��+�+~���F�>=hf���F'o����k~�{ҋ�E��:/�ݏ�=�	�8�8g	�5m��5T�^�(�gP���DVn�x��yu���Kx��6錓eу�:>3�W��5zS�d.�������d�6A��6?n=yC��AZ���Y�M,�$���vh�փZ/_tC]�G��;Ҏ���L,�9�Fc2"��W�Q��=�3��]��uG$M���t����H�.�h�z�9���쥲�Q���Jkvt�5J>wF��x]<�E���p×�F��޻����g���ʪ�,���:Q��3�L�G;��	�{/��u�z��kT�O��!��������R�~Ee��ƍ0��=�{!n���iV_{�`�f��=U���F�	"����]͙ڹGM�b�:�N�E�§��U]Z5{�x�i��_��V���f܊�J<[0���H��{�ۂ��z���Ջ�P������*����T۳<��D�'��X/�E^�~�[�U?
�ڳ�b8��:3l7)�T͝��'� ��*���"gi�)���1��)]�zQ����D7�O�2��p��Sid]����j�Y��ͅ���HxT=�Yjf}��5e׭���釬��7�4Z��鐆�!n�4Zv�gk�
�a{l��
k�
���ު,\_�����FfI,�R(�ق�b�0��i�3{E�I�{��i�l��r��c�)U��E�����Z,H^F�d�sԡb��<,^=F��f�3�,�*i���!�Q�Y_m���P���v�/k
�ヘ�!��p�ߍs�<k�{��~)w$�	�Ɗ�[����Ϩ�ѡBm�-��E��j�m��Hp��K<������8��E
��G:�P�77p°��W�s�!`;���fT���mG�����mǵo{_ņ���0{\g�fi��L+F�R:w�{ٳ�!f��Ip�;�)���8[�+�mvhֻsg��	�_N���a�%H��L�C/��3,�����B6��rq�{tFex�n��X�ч�����<0�o���f��u.,Y��0�!���f{z�}e�vHf����ah�F��[2"�U�{�[��a��!��/���0��%�d�*/�Iv��>�;]z4�37Qex�N�`���f*�}Tx~4jݧ)x��Pz9�8�5Gi���B�,�5��ŭ�!#P�f���������"�VT0�F�Q���aeٚL�U8�;��Y�f�a��â���B5�����j���!����"�,�fj�Y��.0���k���vQ��0��E���e8Yڬ�wB"�y�v{�␏wWVa�ʆ���Y�L1��3�3+�D<f���}���5��30�6"�f}Ų�K��D�|a��Z�TY&膰��b&a�N�22�/�a�Y��a�L2�4��+�����E�fð�٘f7�p�y�G�6y�fف]4��R���.�0�z��Ғ�F�ޮ�z���0l�H���/	��S�
��"�G�R�C%�"���
yy�P���}�G펞��u^�ћ�8!z�̧����<u��DBy���w��������{L*����,,���4���'��Y��+��c�Y�
<��K"<R�i�y�Dn(n�\x��!ˢ��
Dͽ�8d��7-�BͅU��s�/��]p�����s{�4XC]d7T5��:�H[�S�d/���e����9�*N�S��j��)6B��o�5�;YxQ�E5�4��G��Jv���-�����C6A�^>�ѐg�s�ec&�xc�Lx1�D/�tu�]6R��a��MccΌ�̄����!`Όt�yHlc3����c83C���١�ծf�A�d7sd83C-%�Q�}'�w��~Ă|�ᒐe��d�c83c0f�K��³�>	��by����I����V�C�s9تUR�5�T9~.��F��Oc�+��=0��"lZgN�����}Stܫc��6���}74æ��[�t��h;��b�g��֭����L���'"�"��Z���jҜ���+u��ڰ��Tڵ�f����i����M��I�k�,z�)�wU��wO8[V�V����f���5�Sl�M5Ӷ�z���p��Z�8�k2#MV�y�m]�/Zƍ��>�4r�in��4�pcj&l�����HW�'��J���oc+��
�%5������C���)��j����kT亭���6`�6�34D�uǮ��h�s�K�J����U�؜z��X+y5{�{~���Xk;=���ȿ��V���7�gL�ǵ٦kf��y;T!���b�s^i�ҋR��z��.Պ�λ
�Ͻ�Y�fQլ��k7w	�'e�����ۦ���;�*{��8�a�K��:�Y�Z��e7�5�є^���G�QO��sx�z�Ƴ,UJ�
V�+Y��[�{_&M�rL��:;n�1e^��zuVB�>�[���a���qp�(͹��Y��E��8��S��ޤ��?��'��������n$���p���&'�X�?۟���"~�l=s���ˇ䞗z������k�|=_lBz���q���zܟ!�'�QF�m�Ѿ�jk��^)-��׫�3=�rq;M���mN�����m��q8�N'���~��O9$S����q8�N'���q<�ȜN'���dN'�����ݑwwIrq8�N'���q8�N'��Q8�N'��{kw}rq8�N'���q8�N'���"�Nvt�ݩ��qff8�N'���q8�N'���q8�N'���<�؜N'���q8��.��"�N'���q8�N'���q8�V�{��wb���[��u4�i��q8�N'�������x�i�q8�Nw^��jq8�N'�31��q8�N'^����?)&ɱ>O�{����w��wb��^�ܜN'�����M����q8���7W��w�_��ݿߗ��n�W�'��x�i��q8�M	%�����R�.�]�E�9/dؤN'��ӹ8��)2{��D�̘�]����r�y�)˹8�N'��E��$]���q8�N'���q8�N'���q8�N'���q8�-�D�q4�(����绻���3dq8���1��M����q8��������[��qn���Rq�qlR'���qL���yo'�v�L���bm4�q<��弟'$�c��^�{�[��q8�N'���q8%��Eɿy��w��������b��򟓉��s-ww-��Ir��8�N'��ssw�t]��D�K�8�N'���N'7wwu8�N'���q8�N'���q8�N'���s�H�����8�N'���q8�N'���q8�N'���q8�N'���q8�N'���q8�NwIrs�H�����q8�N'���q8�N'���q8�N'���q8�N'�����{�������x�2z��	e�q��`�c��87%t�e���m��m�Sm��4 ��D�1L ��8��D�(����c��D�(�(�L'�0��0$q�D!8���HB0�B�)D�){<��Fa1$pB!!B �\$)Nbބa�! ��8�&1�,2bA)	b�����5'�������s�F��ԉ��q8�N$�N'���q8�N'���s�����q8��]�˹n���q8�N'�J!e��"�/�R(��J0���9� �!	�Iθ���) 4y�טB�$�җ�4����܂$L��a+B^����A�QY�*8�����F��v���۽
'"F8���m��ݣ�"����^����U���wEUz��"˚	�nD�$K1еR%��;��Z�ƽz5���v��Ƌb1f�^j�Q���Y�]&I�.]�w&�[[	����3mWg���{�m���eW���9��L#���gs�*m�ݭ��ݺ�U���R�-9SQ��Q������>t����q8�N'���q8�N'���r���Irq8�N'���q8�TN'���q8�N'�Ē]�E��$]���q8�N'����'���q8�^���N'���r�O�����M����q8�fdN,��[���q8�N'���q8�N,�����q8�N'����y{�rq8�O32wIwtI%9��=�W�E�_ו�Y[�˶����ZLMK�6t��"�6˭�I���4�F7����]Y{�*n�P�Y6�$WgAŵd���6�^}ݝƲt�M���qۘ����F�ur��W)$���Y��F#+o��i4�9$]���q?���qf�j�Nw~�w'^���"bm4�q8�owu8�N'���q8�N,��[���q8�N&&�M�/wGߝσ�������y^AF�3%yd�V��㼮p��&�G�������9�-�D�q8����q8�;������e�8�z�r�%��Ua!�������K���eڅ�2�:˖��a��%S1�{U��(��Kk������O��p�M��c���v��m�-��I�M�������XL:H;mdp�q��������r"�&8�8H�/q	�!�b80b N#��@� �G����B'��0�F0d�B���
Qc@DR�Q� �$�:�0P������p�BBp�!7�1L%HP�^�"q�$�pb��	�c��`���#D�ND���&(��S�1cB$0�� S0�1>���<!�ąD��
$���acT�R�2@sһ3f��a�y;˵NN��yz'���w�w'+���ܜN<m��^��]���q8�N{�ܻ�rq9�P�Q��v���J�%B��\Un.�v�m��Uw2��Y����Gr��-7���6Xq�I�"���۪�W<vV��Kv�m�p썸�!Kbd�휀�T��j�9�D�q8�W��弟';����H�����q8�N'�����{{��bq8�N'����{��q8�N'�N'���ԓ������'9�[��fb���[��A<��qt��8�C���pN]�ݧ��)$�E�޸���-�����I˻^�y��"q'<��:�N'n��p���Z��E�vL�n�w�8۷CSmfj�ڻwt�-�[���'gnT΃�M,F-���̔���$�FMA/j�]��MbADڹl���^˳�粪��z��.{�w�%6
滝��Z�h���iz[��7v�T�N������ʌ�T���3���98�N'���q9��r�]��E��$]��绽˹w'���q8�l�'��w�$RwIr{{��bq8�N'�����M����q9'ݴb����RX%UJ�29�bU�>��|���_�V*땨��׵��{����T��d![���o�竢q8������b�8�N'���ZoZ؟'���T_+I`�˱��e�wy��������:I"��.��q8�N'���q8�N'���O�՟V���-i�IZ��H;��>B�
+,r��9>N':��D�)���H&0�Q �1�;(��hR��� ���<1
aH�)a�iꐣ4UL*�6����r�"c�)�*nMqA9��E�D�$e;s�|v��� ����:y;��\I����A#ęn	���[���YU�U{�Y�,�m���vp8L"��NwmM�a d���S��J.1xC�{�.>n<KO�:�Z�kV�7V�h��a���aG	��۸�/%��S��ș��%'u(�a�"BC{�q�C( ���BdK��Ł d������"���oV{��XY��w-UU�X�ڷv�`H��a����wHM�^��sNM�Ф
Cn��H(d�jB^JMȽ]�1ob��Db�E����7����������^R1���y8�$=�)���8��L���e�aQqa81�Lc`̈́ �J&7`KD�n��� QiDCKaԚ�JB�؝�T�1]��$�LA�#�a!�m��!!S��҈�*A`|��R=j3���D�R��|��Ԟ
t��j�u���$ƃ��\M���j�:]t�,���nq5!�o1���v���y�]:fB�Id��d���RJ�v�4HNz��b���I�{*V�{���=u�n�,��S��GlQ�^4�%�.	1���b��<��!���'B��R�n�(8�.���(�Sq2R�)L<�^�<���i�Y��+�Ԃ�k\�0źI���ѻ�9��=:��GuV�D�m�ԶH��,3��W������FDڢGir�lu���89�qck���U��l+��ۇ�1�gv�����v�{��ns����3��^Ju::Ŝ�s���:��(��W����S���HΦ2fvĒTɲ �ۇ��Ms���C�1�D�/Zv�0a0�HAt�(�1
'b�!B���1�L`��a8���'0�)��q��F(��H'$10S0ZQ(�Jc�)DHcrS�0��D0C �1S��JC��%(�HC��b81�0�La=�b1JPJb��%!D� �<�	��K�`�� QaDkԟ�g�����ٌN��=v�g�UE@b{z�����r��G^7ڢ�E�����G���=f���>���߯�Ro�����g����5�g����� bu�0��}~�w������^�z>o��~��/F���</��q�>�n�p�̢�1^�cUc<3�>��kh�x�M�f]�ChV.��9�ȿQ
-��5�<�r5�ӼY+���0L���XC�oYTBE�b�r�Y��2�J�.��q��4����xs��ݗF0���Xm3;�{��i6�?=m%����L�
:�S�Zx��u��J �<��u������p3��x�ι�ߚ�!����� ���b��h�A�Ţ��0f)�,~81�];�!2n��]��w7
�9�|�j3�j��x�=�Q��r��Ǉ�6ZL83^�4��cE���m����6?߆-�27t`čX���{=����G1 ��� �V���rv3Ύg��1�m�Q)�+)����7�x�<i��qRX1�FaJ8O�����qS7�^�W�A#����V�W�o�G�cg^|��6E����� Z�Y�n�gG�
0Vx��OZR��F��k�E��������$��e�+�Qb@J�DM� =�T7.�c��:mS1l5u�u���5��]���8�`c�����cFش��	�C�R(����/w��)���)�A��:�4���y����4��Sd�"n"4@�d@�G�%E�a�Au�f���G�2�U�����=��u^�Pvn�x\�;L�ض���8�CO"�8^kq��<lI#�7���R{�V�@yVa�1}���P����������#`���s�}��5g#Y�V�b4��WWҼx���=o���e�����2}�{��qFb=��b�kfaE{��_��b�e����aT2�~���>�~��<a���m�n8�x�iE�L	FPU
�˧��=B8+���:�Hy�c�F�5D#��N8�?�����+��o}W���CM��7�n�"�;�H�$�Ѥn3Yܰ���ǎ�B�(�e��e����~#� �8�L���|����6p�)��ߙ��u�����ǉ�e�<)s�#/���uS�ie����<`��B߉E�W�����ӥ��#
��:-/y�g�h��}Q捳�c痚�߶E���5��s��SE�[��A�v�<z��Q�g�<f�4�
0h�g�0k��Is������!�p�i�k�����h0bƫE�íh��5�{�\�z�ෙ��P��g�<j�Əw3����p�����i���EɌ(�Aɲ�4G���!�h#IYǬ����ߌ;����/�E3>�Að��`;��x��H
�A��=<?t�}s�����<��GY�� FaXs'�p�ޝ�42h�exK�Xt]�s���9���N-��F�GL4����V{����f�9aP�7��zY�d�kG����M�����h�6n��"�=4��!b���E��g}Y��٭x�kj������G��=��єc=e�_O��gq[����2�+�A�Ԭ�����_�S�-<x�8G�U4,'�qF�"�D,�Mt�g6k�	�ᡧޞ;�|�4�3rix�i�eX���Cŕ೉C8F�;L.C���]C�Ǿ��h�x�7�������-��B������{�.��v�W�K+�N��B��q��m��9��9��)p�� Ѝ���ǅgX��qM�x�e5�3�b)Q�
�a�-��\,ҋ'x���#�3��<. ���{}�=������E����F��h�N���0�x�,ê�� �����h��e�Qe���YDVJ���3A�D�W�M+�=�G�M�q��"�����Z�_���H����df=�eҴL&T�U�7��vi�aOYl�6�����#F!X0�,�S<A��'�k��Э�4_4{ƖQW�~h���ލ�t�̧'n�̄i�?�p����a�r٧�V-$0���*���/7c�~����_�1駝zk*�3O"jͤQr����m��H����4��e��6�v�12����iE���vp��.N��^��Y>���şY�N1i/�)���e ���A�����ՖKf�a�����Yʸ���L<av�~3�=^�g$qP0��}�d�f��4�tzy��Q
�\g:�̦"�E�/�Yc,�N)�8{�S���}vW��˻�z1n�x�b����}��%e�c����o�O�X���Y)R(���H�}F�{��B��q��i�Fc���1�l��N�ͱ��7��p��:�/�3V��FU:��Q��=�Fxg^���
���ᦡiC48E�94z���^�3qæ���e�mx�FuK��z�qd鳚#42o~=	�ǭH��u�F�T���~0�?Z;쿽vc���T�nw�d��1tb�/��J���cåv��{�%�vB�us�!�8��*�4ua�!���=�1b[E�4_h�Kw�E=(�Q��<xG}{�Mu��JR8(��E�t'����҇�yjv!����X�J�c��i�s���$� �������θ���<z�5B�BM���� ���|����φ+38Y�+�r𫻲� ��o���y׻K�r���Ĳ��
��k�k:�K�ɢ�s�!����Gi+yǧ���70�+����ֹ�57���#�J�.�[�����k��fw�Se�̶Yk�%���+�]��3��D�{��l�P��ɤ٬N�F}�x���������TBu����Eݩ�<���}b�f[Κ.ބ�����0c��۽!`ƼU|�8C�x�?��(z�<`��x�|��"|3�|{�I�0�[ӫ�3��c7�f[��E�o��j�;��|`�_o����M���Ϭ\b�+�FqC�a����2隻�k4��Y~4��CRj�au�f��<t���]U}T:��w�����{x�lk��j6�Yb�zh�^������F_ЅfQ��y�0
Y�F��5���׶D�C�f�C���"�0���"1	 �����%p{&����t}����Ԩ?��Y�Ɇ�[M���3�)��X#�IZ � �F�l�$E1Z�&"*L`��W*�S�\i&��ƶ^��  2 (������tnr�k�1
	�BX�@l ���6��GuyL!���0���1�q�a1�@��J��"Q(Jv�${q�9+��a
@��+F�����cF���q�����ػ��oc�ȏ�v\mfn��˶�)Y���v��N�#�.�ܪ��<�z�{�s��5���U�dv�QXVb�3�T�\��݄k���ocBA	��0��ƌ"$!��#�&"=���� B�Sc�o�6C-�l+ˑ��}�I�T�=�/t�U�U��w%�+Nz̐�ܫ��n�7{��kiG��n۹�v���S���c�]I���N���p׎"#���E>����!9��=�"�HBH��6̻v
a0��1�!w���&Tk{���c��#��q��"ExL�{ɱ�$'�u!3\KWU�	�R5k��fm�,�WBd���b�q�8u�t獭Ӹ�Zq۵sF���w3smڣ����U�]��M&�gRS��aH�1�z#"#OCJQ1HQ�B��B�a�0e7x*.$C��0���O��1B�Q��)�Ņ���x��\����gJk[�oGa�T]�!s�.���k�R�&�eH�r���<TT"e.���ѣK��+mthqh�[/R�.7
Ҍ<_ѸqE*��/�3����$Z.�a�`q�)�a���T����<a��������(E�C�r��,ҋ�gҾb��+<�/U��O���������7���l�Ӆe(��B�G�݅�H۰g�4����f�Na o����)v^*9��mk浵��S~2k0ᔨ����5U��er�gj���!�70h{G�|��D�Y�9\���:=L$+H1���m��CkKEs��Ni8��#"�M��nW'Ny%��ݻ�W��9�ca�&L@MȌ
j�شLRR�],�J��Bי�IӒ��C�F��h�ʍJ>��(��,e[��� hjE�(��H��c;�i�O�P<J�!!	��zg�Ri4�5aM$�zW�aa"�Q���z��c*1�=�R���=�� 0�k}礍��ߥ�Oy���x6�h�m��yS"��`IA(�9!<�=��v�c�q �\�rҒ��j�&p��}d1F��� �8���
$���#A��[@T�;���9�IA0����D����7�oֲK�]�Ff��	�Lp��ӯ^TԖ����!B���F������(oi�x�H=Y�e���&��|5h�80��5~���Ł����u�ޤ�""a�-1iC�+��Ȉf���=2�f9s@�[�K��~&���P��,����$�h£Hbئ	�=�Chiш�#���zҌTuv=�aJ�p��;��Z�ws5a�n�^�ٛWܞ��*�FM[�fĘlt��1���v8������oP�7��<�s�������q�ɛp�R%�_�u��s4��$���������Ѐ�C[����b���w��(>ot���C��^Q�145�n�{����P�w��¹�ۆlbخh��Iǩ�fZՙ����|��k$�-_�6��I6����g��F!#��ip��NG&򷲽z}E1%�e��I�{j8����)�4���1�N�W[)fb�a`�{ɽ���q����1c�О���ܢA��'Y��۞izX��C�y��U]��s��� M��H����m`���{��0���X-��{�Vi��4l�},=q�ykΪ��*h|(���:rQר�J0�R0dI�F`�1nl*�gsªF����|6��P�2D���5؈��o(4f�6����j�@؞�����j�u�A�}rۜ���#d(�I:D����(�"xV�2�`�n�zG0��
oz�����E���B���D9G))F�ϴ�TC��o׷�4bh�;�G��r�1o'�|�R���hH����7kG�RYIJ��6�lU��#FѣtT�D_5�h�蟯�D~�x�߮%�X��_��B�B�2(�֚ͪ��̌휧U�u��X��iUbhQ;��8��q"b��z���ݣ����»G�)b):�`����	�7BHƙ�*"hޑ�[9�`��F��o/�	��/r��6'�|��{^#b�]�}�ݮ�Zj�f�� <�w��Y�e��Yuf��
A�HLo3줼Z�<s��ث���F��ŹuD���l&M�8����Si��6F<�M׈Caӱ)���[��aLSSdHcv�z6���O5��L�DR��*��T�Iܓ�C��)�)�F8I�C.^��8�/$�������}����n���zn�w�״�����lN���z���r�Z���-�Oy�&ڻ�H�n�cj;��u��p�ѭ��wځF����J�,t��f�e4�fF�J�������X���f軟c�"��-�H�sޚ��������k�Vܺ�$�>Pz�����B%Ϋ�J�\SG1����7��t�g�`B&� ��i}w͙0L0u����ܓ����KL��x��cc0g��U�C�AF���Y���A��wf�ď��~6C���b��ގ�(���>w+���2�0�}���iU頏}�]~��4�D�nii���HW�>��}SL|�s�=;�y2��iǫ�y���O!Gz�J�T,�z?�:2�xLʢ2��:����F���i�г��ͮ�����xպ����7���nC�{��3�_��~�.7"��Y��]����+V�~�{����P飡�3Z���>�fh��jO�����(�W�O��K6������5��,�~/u=�:�2ѵgf8�� ��Dp������\���L=�����Ȳ�1�z~>G9��3_0ֺ�v���Z~�Ό���B��&#K�g����A�4h�S�C�"���0�O�fq�yxr�ǧ&�p�0��C$#�h�g��iy{&�? K
XRIaCl3�kZ�kZۻi�gK��p ��u��B7aB�wN�����sZ���[d�!	$!B��~fL�!�L�{�pε�kgf�#7E;�.�kV��r�;.�l�Nk+�ܹ�{�w=��[;g��Z�r�Nk�k���[aBw��j���ë���/�V��*�λ��u����{����l|{p�<Y_��xgQ<Pa��VEHEl�9�$|{�0���`Cg��^&�ۄ69\;��(l�i�<a�Q�/E�f�����Y�64SA���4f��d��U�����E��i�k6�Q���x�4�>h��h�uk�5:0�čr�;3fXx�1�h�w"��p�-4%���5�F�t������Fx�f��iw���f,��P��%X�"�Ibu��3��8h5d͕O]������D�-��M=C"�B���=D��u;���"OD��zg�鐤�cN)��j/R�H��g��5L(m.}���am�%�؊��05���9>Q'y(n�B��4��u2N�ipLEi`D��E�jM%q!,�[� ;�i �{�̤p�w,`���r�՜ńr�,���0}b�DUWֳ��p¡�mVA��Eu̲�/ �
؁�1��,��������	�t��[�	n!��z�^!��Q#�^����_��ic;���Ϙ��&� ���	:����a�d��	8z���n	���pn�ݗ�F%�
rQv0K��f�|L�%�m"��A�X���r¦�]�B⡸�`��1.�H�0��0-P�TM�D�X��c��U�U�# j*���"g{��@:pc� wt����6َ+6�I��Jc��n��I+:�,��l-�
,�q�w��y�g�L%1��y�{�U�,�֖�/)���Gb�..��&u�b���*bdh�m�!��*n4�|E�"A� c�/��Bz?�$���������H���TR1�L}~!cP�����i:�����1?��̃��$E�AE��`�9޳�0f�a"&��"��\�r��f$0��r�Ca��S��M6�i�ƌ�{�J��1.6��?��L�)�ش�4ig7V�j!��.� XSqJR�(ɤ��i��⓼���� ��sY���6>�B��gѦ��+$pc?�|aY��%+	<#�h�K>���rҜ��P�w�E�>r撌1���qHy1̏-(/�'�����fZݾ�CJ4��&��=A���;�h��B`Jc]LU���`Ө!����z�E.9͚��XD��#�	��pn��s%�(0��l":��߾%��4�H(�
O�v!@p،mAօn�oBi���"�@Q60E�D�y����5�`��4���I�9_�J��<=��ᄆdz��	�f`���#���u:������h"��c�y*@�#Ak��:H��C��W�H���w2]�.#���c)0�1�J[�	p�O����������n���̕L�-o-�!��fRǎ@q�QR0"�ʛ��k�����Ȓ	�H@�y �k:�8&B��y ߔOQI�,����CK�\��g+��0k��I�6n,,HAe4�&)DH��40�F���E�^�TN'(��v�MB1N���pt���� "��� n(��	u�(⃉h9�;�$�p�P�m �s7�2�tZ[��D�D:���������� ��d= j*��!����j,�kc����cg���+���d$$scۻ�=���Y"0���>oǾ=qbu�fL�+�M�$d��U0��f��Ƃ&�.&a7S���5ڢR���j��i�D�)��
	u�'���e?��C��,C�N�-U�z�Ev�;�4�R'T!hP���@�M.4��zZhhl+��.�r�]�s��JH���ľ��̥�����	qV��Y�� b14�}=���c�eT5 (`��"gz޲��c1��zXJ�ZJ$6�0�S�CHQ����(����b&�i;�39��̎�6�}��\qC�Z�H�`6���RU�0A�60��F�K�,	72���y���(,3������(�G� 3k8Rs��+	B ]`��L��~q��W���� ��+�g{��"u�'X��E
$t�u���!d)lH`�&�fS��W�"	P��{� 3J�zW�QqA!J� ��"@��)��5	��<˄��������ߐ�sA0S�@���!e�Ó"$H�H�9�3``5IAp ��D���n"�T��@��4hk�D��:�ᒖJ�Ŭ����cIy�хg�Ś����*Hc	tLCT*U�@������H/+����3��a���20\D�aP#�5|�@�-+�R��n@���I����A6	�pM#��!pi�߶�rff;%�.G/r��fmT�5]�Of���Z�k'��G��4�!����mUx��c���ܒ8��%�4���Ԑ�ߨ�]$������P=���Ϻ�aE�|�Q�B�51B�6!wzF�
D�E�Cb)� 瓖��(n@�E0$�� X�U�]��)bi �8@H&�"@;��2��c��!��i"�� �P`�^w��U���Q(b�n*=c�J�9w*�.*��*����v��:E�d����^���L��>�k)���ν��$c���ӹ�\3�[����~M����L/I���_d���ѥ�g��`��S��4�U����0hm��ƣ�F�����2195�9��q-3�6�5�A��s�4��M�nh{j��&5G��q�d� �:>�!���͵��U����0�5Q�5�����Z4y���G�B�Mi��c�T:B�~Ӟ��b_?�a��0����:Q�CшlK$M�8��c#1��)���z��i����2̲d4������M�|<56<���0���;xrVk�ŭ�F�?��L:r��9���/���y�<B��K?A{���U�[���j�w����?��g(��O�Z7$����担=�?�Ѣ�vU�͜�Q�'��kG��͟a�,ŝ:t�!�Bg���O��'��JK�����b�D�`��>�y�i���I�^���z'��hafH���i���l:��U�Ø1�'TR�B���		��Mp�����s�����z�ǒK�)W�����u;��T��ms��ʱkm���ݭwf�ꪮꪹP�tܝ����H�8�Bla1�& ��1Lb�/a!�.ͫk�B8�8f=��E�ȳ닺�=�d)Ysӭgx{G{��ݡ9p�>q�Q��/��슭[f�7v���;��h��l��Y����)t�ݴ����HEpJB�Gov-�d���l�3��c��O���<�!
A7�B��0�H	LA `�	����%�-�$��.�Y�8��5�%p�tf1�tKe�㌻���gE�Xɯm*a#���2ɜ��.ee��](˗�����S��|$v�xv�ӫ���1	��(��
^���/JQL"Bv)��ӝ͵�s��(���qy��e�u�"	��"\Y��<:��mt�.&$�F�hB�t����v�CL␤�%J^��9
Sz)8z�IfYmF�siiq+��8Ŏ��B�Y'B��HG��xc^��wN�s�u$g;��va^�[7lvΕN��:ҝ���"A�	���'���H�c�a &)�c�B�
_�{<�ǻ�����B5ۙ�]�50$lj�7�Ii�7�Đ�!� �І�awʍ.'��-���&n�(3!��h^�G�����~�,�<j.��L/2��(`e;�L����N�6a�T��48e:A�8q���3�3b�����4�c�k)�]iB��2�V��)n,޼sY���U���1x��\���NA��XCf�o��t�� �WMgf��֩Zc��C(�X�)774C�4jœD��[�g)a�~�����ӷ�g��Щmͭ��m�@���2F�O��ٚ���<>�*�Ȕ���	���B��MrV{[whS�����8f�R��
c�7�bF0�!%0�k.]І1�,���&���Q��)�K�O�?��$��!ܔrm4�Ψ&E.TȦUE"�
2�F0b4�z���H+��'R�Pys������i�.(�P��T���H-$��|�j�	7���܌\Do��T�(S@�61j-$X,4�9�sY����`};�a/�1ۛ[��is[��s�QK*��'s96��&�;�AF��-�St�H{��zn�qOb"c��1���;�`�1D*����y����7��6���b�$�p^ӕi��&Wqr0�n9���!��盒O?��� �iq;y�{�o�LB�$��$刔����(�hN'!�w���x���"�Y�����]��icA�^��Z\CM}�8� y ���� d`Vs�չ�hzH�pt1|��T2���\h�9>nH���J��'�y�m��OD�E�v�NHe��KH��ttG��A߈�"���7�1���#��R.�`7(�w�yfsIA�%.��SM�[�]_.-�pm��V���+{�י�2�Ynd��͍]ͪҚ�kkU�*�j6�2�ҁ�QE'� �؎�)�T�-�&�A�4�?}!I��-7���/1�F��ʛ�(>@Me%!��v$Ђ0�ۋ�и&`q��F!����Q�CZ	��7 o�g�f���BǨ!c2A�./}�<�JL����A�\�Z�p��ZcI�.��	1��ҝ��0ib�{��'�'�R�*nQ���RZ
��L���-�]ٓD�Uv���;$F�=�XF"np������͒�v�����GAC��y"V7,"^��d:!&6�8D�ۘ&8���f��:� c�sD�V�ܣ��7$/V��
7�G��c�!�Z�*a�4��Ithq9X���!m�����D�qo��\Ն$ �E��C#����\%��\A�@������f�2�/0s�1�NZ�_ψ!�;����F�"9��:���Ƽ$1eB�R����.R.�`��&뚙 dM�x�@�0	"�/fΠ6����Q���:�F���¬ ��.�!��\;��`0�`�����W��W�^e$bR�0i�sS
���lZl\in����8��L�#iH%ݡ�!?�6���%�4�K�01�"s>fƩ<������t�yߛ���X�b�=n��Ǩ=$^N�+#�d|��0��E�Y;�`5�#�O��HWl������iq�o|�&��0���DȲK2LP��B�#���i.4�b�"��r����7PCc�_w��r����Q61q��3�di,]�]A���T/���B,+"`� b� ӖR���L6�l���F�2K5�}��#��u���*�@�h]l]�c�s�m�;�� �[���<�c�a'f\�!:��̥���q/GiP�������F&S��b�.������<�p`2��72]���}떘��f�1-w)rH�.��\99�ȸ��W+�ך� �1q�[���~�?Fq	6Q��a#�Hb	��d�!M2^#4ËJ��ĖA�MH��n�!
B�)��6��VG-�\�b��Ytф4�2Գ�B��S,h�*���`�p�����J��!���b�\Oa=�!4��{3�������6�j* 4y/���+����1\�RS����H�9�s#T
MȐqq)��3���E۹d�"��i���gAN`�Ļ=�H;~�e�6-1q[�&�S'ŋ���&�vHULN[m�TY�A��Z�#wʙNPPD��x���4�$Zt0�!Ԩk��ZD�@��L�v0n7�����8p)&�F�F�8�k~�E����4{�L�I�7+�b�b�i�k{�B0�[��$�'P�bu�פx�0�F�#�����`�i�sf�.(2;HB!��"D�3ɛjW)�e7�H�5��>y�����/�U+=��Z�;^s��ߏʇ^54���G}4a�S���1�vOC��B���3���<n|Y����Ֆ`�&��>�������?T��R���SgiGJ�ω+,���JW�3gxhᆾn3���R߱B����n��ꆚ1��[0��o���Uy�x�:Y^7�~����=G[�xy�~'O�o�a���Z �!1Zx��4l��î��`�o_M�/���=�ニ��F�]t,�q�8e��E����"��Ær0�~4���ʅ}T:4s��=�&���)���#7�Tvv��}�U�a/�a��3�=n�BB�!I#��kZ�kZɎsGN�]��V��Jʺ.�V�Zִ;��]Ļ;:�WY�r�V��c%�#d!B���!B"򕶫U�kZիZ�;���ZѭZ�:�ڛV-XsF�2@�(�(�d��(YR����k]6)�\��̖��5�{������>�n�K�P?"�d&p���Eگ��Z�V��c���Mo���uT+��R�c)�t���r�L�}����w��0{��/4�������z1Q�oK6��{4���X3�6P��eP7I�NR�ʦ���f�\cCE1k��6�6`3�Ü6f�#���g&�Nl���$�����Xlֵh�k��`�����;�������k���x�=�G��C��E�2��=�tc2�x`a�[R���&�͗��bx`���E�HB����ya e�E�.v�����۴�-1���9���Z�xSaK�܊�:�V
,����"PA��%Ev�n�|�����60J���\NVi�L����;H:$`���ª`��U��#��^��e�����0]�ֻ"M%�]b;f.��3Hͫk!1�����t>��C9��C����M/Oz;���d��Ɔ#_!����Y�P�FKa#�&F$؆�B�zp�<�׀����$H�sY�2P`- P��i ����r�6�7�.�)q1f9��$��i�{Q����FF��4��������>�X&�is\��B;�p�2�d��m6�`Lar�����;hBª���s-w6��;т!0q=d�w\��PF���݃ukd�G����	{�������eF9/f9�R��2��Ҕ�����"c	�b��=<�p�U�x$Ix�b����Iڄ�Ǽ�+������9��9�4;�4ad�P{�59����"�I��܉��<�� R� h"�.	����4�4#�O��r}+n_#iF.4-��Ñ����9L������a�a�"f�=8�D��.R.�s���l�bR`0ġ�M������4wT�c��^�/Py����L�����pz���D3"G�#QC]}��>�`�&�)]��.��0!�~��~d�&XC�HAy'S��$�8ݴ�9�4��hM,�-H{'z�d�d�r�w���%w��@�xb��c��k(�m�u�������b����ipLF1O���Ub|>􅲳�m�1q����N)4h�dY^	(ʻB�z�gZ6�HN�+�@�j�K�ȝ���1�I`H��bܒNA��nF�#��j����b�L�0�F-�Ə�!-S��9,��Lw%��s��ݳ6��ַSvi��˃�d�O�����}�4k~ﵕ����=�r����σiV.	�Z����s�B�	u4�NfHP��l�-�	v� e�ԁ7�E;�|��G	��k�L��0K��;�FƘ�]Ĩ��p{�'y����6�J���qo�㚰Ʉh!�џ|���p�"����4�w\�mٽ܅e�,v�3��蓄؄��DG>z9xϣ�����or�6��,��TvcLa��Hͫ�ٗM'Df�� ،ө��z���T�C�"8�]2b�H]���Iw��+���N������3�����r��jK��$0hQE���wQ����C �^@1a�����`(���q.@��{�3t�d,w-"�.�/\�NRXD�7#pm�Ǝ�^��E4�O�󰒿����K�D�n&��f#0鄦�-��Ͳvt"�JmaLU!�'2��f lb�K�����@�@��#�P���8b��yF��7"E�.������%+������O+>X�cK���;�1{�7sxi��0\CK�|����G+��"��9��~����Am=�I�@�d0���
�P�q��i.1-�.����2W9V@�\���@��7�w��!����C�9H> /O�{p�ց�����2"LZ� 6x-��Ǚ��
�#LK^�����~t��|��4�,7̍����w$�a�!a ���S{�3A��iV��ō��y�ٿ�b8���/��8-61&��"�7�3uan�;�����&�����Uu�uWwQw:fҙ�n�e��31ܥ���nd�Ѩ��w����X��LX�w�8Lv7#|�C]><���a_���PZ����]Ѕ6��B�7xw�lb�"�c�ZS]���Źq;�'3̅�2�)�����g��	abj&���Ŷ��]{�	�6�T\l��cF���_���@q,�4�����k���<WEl��{�x��'5��Æ�6p�ï���~Tv~8����*�~�3�?"�B����O���_to����xL�<6z�����Y��h���E}�z/���C&�<6lz{1"���)��L��61�X�ҟi��`Q�3���ސ�ĺ{m�Cí":Ņ��R�+��~\M/�+TFд0PbTh�4)G�!����n��n��n�f�X���{
:��g��x���N6�U�?q-���}.���J��~�4ɱ���藸z�xdk��t|f��Rd������1�5�'�4�oܶ��(=_��#�l��j�}�ǚ��5��O���/���v~9��/zx���8�(_L+�ip����1ҭ�z]�џ��Ӎ��ٺ�^�Z���ڸ��Z[Eڻ�SN^�V�j�U�ꪺ�UN��ѓ�zLb ����1"&)B�l�c�0�`��I�ХDآm�vɉ/e$��|��ɷ���8e��qs=���u��[j�i]5���=�U�����q'ik���m��E�v�n�m�&y���kʈ�mn���厌빤�^Y�\\&*R�DLA1��"y!1�0Db8� }�0P����B�b�È�g�"�fI��E�5�M���]�չ�V���m�H�#�n�Xl0�mkέ����3�EN؟]��歺ls�.w�qp�1�]\E���zݸ�ɌG����G�p�q����a�h�-2�ZIF�YyG�q�L�ܛ�}nc!�P�.���Rq�p�0�	yi�V�q�cM"D�q�"��bd���F���a�蘶D�3-��ͷW�=͔yڵ�a��� �1����L�4�ôbJ�@�JM��)[Rh��d�as=I�;�8m�q{�� �SA�1
"$0P�B��1R	
A�
"2w�����E�꼰e���W�T�(�f�b��p�٭ze6h�☻�Z�١�<:3#���뛣&��e	��Ž�j���#F-*��YB!4!.��xE<q�C!ة�چ�\K8C�Q�p֎S�|�A�)��q�А��8p�����f�N��!���!9� VRRP�җf�c�E�ΔѲ�3�:���<�ei���C!b�_��.��"����=��OH��c�ė�@t泒oR[	U�&\�'%(���0���a��k�r�\��wmƋu]�]�BDq����D�l-=;�ڎt���!�؄+�(�z͈Y� BQz�.� A���^������VQ���(��00�=�-�ّ���J27
�A!M�	�A��!����E� A:��^���n�!���S]š�wޫ���V��\��A���'}�Q,-����p�w��D�=sEk�aX.1>z|��+�c� � �08ѻ�sOXjCN1��"�GV"eCHˉ. ���q`#ǝޣ��Pv��"�<��sPF�m'�A8g�`���a�D!�x��0(4A���R�z,K�iF�$��4z�6i*�M�H1nI��*Kh�x~�>L�c�I�9�k��8��*���H�pti���$�5�X^n���yp!���w�H��pN�|�RRD��K�j� �6�K��J�<�3v�������٭�J6�������w���@���$�CPv0b�_}�Qb��o�
�ѷ5�K��F�7>��lt.Љ	�U�8�$f�����u�Gr]A�@��u�s�0�ev�Spl`���3t9L��.����|ޡ��d0U0M�ʚ�_�9ėϳg���v�c`÷j�3����v��[���C$�3?B<�n��X�i��O��K�;�-y�m-6#�Sdդ���$��s�-([�$#��-j�˅a���Iq���ܝYħ��P�A*�p$/��k)N!�N�A�"퐃�g���-.�r$Z�n	����$L�K�izwő�~�m�l`���w�gy����,����b��,�P2ﮍ�+��1Ӆ��F�	�w�ɅG�ل�<s��0�F�#�ϧɵ��݌ƶJ\[o:�A��`��I�M��&�1"V�!K�`�mf�f.]мB�f���˚� ��CJb�ߣ*��oI�X�
\j���<�
NNǸ�c�.�;��2;���K��pK"N���$���bm`���W1i�p�v1.$��sL��!�����9�X�p�h�a�u�jїC-�ȫm�d�Φ�W��C��2�8���ű�u��1�0��i<@N�\0h����h�w�]�K��Vf
K��01��>��Ö9�t7�'+%�f%&0b\a��R}#��h��f��md��t)1!�Upl�HI��*�R��c��CG�=�}@�q�h\Ca��feD��`�i�F-O@p�;ky @��X:�0n6��;Tv�.5ֵ���@���>��_�+����c�0˩y�G���Ӥ!HV���.1(&�7�=9;qp7 G�����HYa����I��sl�&q��ǌ=���b��(��~I�����K
̑<��m��v]3��wYz�[]�s!.v����
"'��������~���k�g��
��"|�4�R&[�%��Gt^L[v5�[:�Z��XPa,6�����^�1�*8�s�/k�?�1�@�5�s�}�Z,D��Gc�X�/�|\�w�|K�;��y,����iBD�5JDp;�2m�
8���8u�|�φ�:md�D�}����=�ݰ�,้�X�z	Ș4Ķ��7\C�h��"&8Kd��;��E4b4�Ԃ@��L��?
	HC���DV����N,����n�m� [�
N���X���p19���g~ٟIQ17�����9��&1w�V����7j"�b�9��7�
�%�F��u�>2c��D1JPݺE�Zlf��"�9�:��0��h)��C0�Avtr�l��<,�oq2��3�*�&n�u��͘�4p��8���8/�{�9�!IH�B��v�t���-Y�;�,(g��+�3�P`P1ѯ�K����0�@�o�J}5�a����p�>�?��X������p�ނ������\�/|�;Dg]м�����8��Q�=�`��Џc��e<S�gޚ)<{�=JO��_�Op�4{�r��끥b�i�;;j<=�����/�)��'�^�٬����YWA��{�mq8�p_�����W��)�W߽�K^+��\;�#,XJDW8���+x?�]/x|O��ο��Sﾜ�h�6hg�2�������ƛ�VJ@�ޜ�'��<oY��l��c�Q���G�!�����_��F}��fe[��Y�������ִ��*�2HQp��g�B����p���N���E{��O����3�=/k��,���Ą<ad0���#8�a�����x;�A�d�h�x[���à�����}�f���>8Ed���Ĳ@���l�])��C��B���aB��%�!-m���Y�\�K�=g[:�0p��!B����nYs�wNn&�3�kZ��Zֵ�km�kZִl�j�:�gZֵ�t�e���WZ�z{�ij�λ���m�2�nl�ܕ�Gf��]ZKF�kI�v�y�������gd�$ɓ&G�|}4�E� z�Æ��v A��I<d4c����%��@��'���F9�Oa��fd4=��T�{-G���i�?O����Z�.�0�KC=0f���ma�S�xo6�B��}�>���/J�$h�o��n/0�_U|2���_aG;#53��Q*G��R�6t�:�Rx�)�0Ú7��4+7�w���G6�if����X���53�	xx���d:�qFj��м)����6���@��r(xxIw4�qX=��{	�[�@��y�ߚ�7m��_�5�ť����(mg#�s�۴ϾW��/9f#���L$
�b��,![��X��4�}﹦Dш��惙����hȆ0�#�f?h����`��8�?�}��rK\Ss%�e��s���jw1ZX�7$�9"����'�w:�s�b����?��K��f��M�i�a�����r���
xjxNK�(C)�^C!I��I���<�X^�����քE8.b9�}�g��R����߷����4�w�G/�2��=�L�<��԰����e�ʈ�@���C�kɎ9����qm���oV��g�p���)HS΅�dk$Y�-��s+:�)K֘G��#Y�c���&;��zHo#;��]��D�/�'��>��p/�<'DI��i�9k�C�Y��$��
{��>���0�a�i���O��(4o�|zg�偠�Q� �/]y�,D#��n��d�W�G�o��Cܘ�td��0M{B4e)+�o�ޥ����9.���������l����·�/��}t�P�m�}�pa�b�h�����hkG7�?�s�v�q������))H�-�7%K���Zb��"���q���L��Q|��"qk>��'�8����thLh�#��ϸ�n�%G�C��k�Gu}��&^q������T��x��[�1���v��Ƀk�x`�0���$F90\����} 0��(�Ŕ���򒘙�����\�H;�3�����.%�}?���DYiD�amu��S=mݮuNu\ȩ{���?2p�D�H|�9�bk�k^7��*"0>�G�Ylc���N��'�{�4��A��^z��Ř�yIHB`��\Fo�����NV��w�ݏ"%�5��P n}��5C��pi�S&����������J�ۚr��sx �@�V�r�\���Z�^��Dn8�mp��9��5���5%��W�f�MM5�1���CD��&��V�6m`�+'7a��@tC�1wb�)cw��"AX�c�"��;'sc���@��B���C栛�	�l�cg?B�&xÑ����w'��"�H��֌#�A�tHE��� 4d�?"�>��H�)���Pki�b�����Q3p�g�'( ���M'}��"�e�>�����Z ���#��bOR���K�1�"h^z��� M�Xo��s`/Mk�R�H�'��D�
Xa�!C�A��J �>����(0�`�̟k�Ѐ¡�sm~�}��A�9=���R��:|�>d��'RK���v��0�d����Ts��s�*՗��%��*:�����a9M&S;��a��l�q��H�D"D �' ��}������\H*��&���y��d-0��~���3#�c<��Z޸�7L�z���2��Y�$6�j$���Civ�ۅK�y��A:EA��iv�w]�-("op�P��z9��,(+	�]��(�@8g�M���c2:[J�!)K����MtkF{�s���A�;~��	��<x�O����5�N����+	L�nh��<���^Hd��!pdU�����(I$���HM(���v��wʘ
0�[L��7�@���Tc��ڗp-�Nb��7�5 3�ٯ�"@c�目J��7�¨�&��H����>{�c�Cw��E"��ÿ���{$(b��~8�b=��Wa,�x������
'�um�ȗd�����������c����d�M?*Z~~?zv��}3���^�E��b��x�/�~�p�O�if�1�ڒ��}��r*��T����Wڮ�����i�����_��4�i�#���i�P͔���4}���}�*�9���Y&\�ٴ?X��U}��
+��^�tp����i�||Du�|�p����W���Yㆻ;��O���y�(Q�����v�����Yk�a���a�a��`W�`����J:pg��>��'u�����ˍ2���H�Ü��(�d��D�q:!Ɠ^�r5˞ߩ8���}FI(��T�wW�����ܼ�Ә{���Ĳ�C�9n���UU�UGޢ���1�)Ld���)D&�D���aJAg6\�@�(;m�'� a+�a��������U�,�Â�t�]����F�T��w6��]�ƍjn�n�ª��O<�sv�˃+���]�X��;RJU�ً���<��XJ�b�&a+)n��u�a�i�5��4��H\A!D�!Hc)��D���!�#����&�	D�R��H��`ۆR�,[Z�ޥn��=XNS��{[���U�U��х��MbA3t��sn�Z�sf�;C���g���m�hꇳ�g��nM��!%D��D��ԡ����fA5��iԒV�'Z����oLb٬�	$���!H^i
B`a	%�v�m�����"Q1�oS/c�)l��#�JR񄒈��13d6�wdв5�󥍺L�Cnk����t0���bh0�15u���/Y�&rڥl����m��, ��	gG<�p�r[�	P�
u)��!!"8�8�z#�"A1L�������w��z�(K�6g���M�3t�A�>�Yvn�X:<%F��uw�iZO�
<�� ��;#
���o[4者T�jFx�UP�����b�viB�Y�#p��(0�8u\!���p7�4��leZ!����c/NR�ÆzMf��
�l����;�&=��I}ʸ�R�ԃ׋�b$n<�? ;��OѢfEc!����g�P�e���n�:3|^[7��oH�g��:R�3�Q���&Y��ag�~�d��b����<��t��?����rb�m�ŋl��R�zJAZ$�)"��LN����fD]v�fd)���)�w=e]VK����e����"SX�>M��.5a#�ѣ��^nN0�V�\r�;��8��<�y�9����DA�S�NDS�@�()D�r
|z|(=O	�^L���Nq�KD�F�o�`���ܮ#AB��kcu'y�M�*�q,{�7��È3�s�P�#|Gg��6��|�ɾ9I&B���)Ƀ![I��A�Sv�	�1ӌ�)��s��ؐ, oG�K"�2��P�~@JR+R �1Bj��)��a��8��ހ�" D��6�+���)������N&��b��?}!I��o�f���)����v�遍 ���a���,��=�h�ל��Ҽg6����a�[�L�<Ult0��aP�<"~$9�DNEN�!�!��Ds�z��üHyC�����D��}$nWcJp_b���
΄Q}��AU��(B�e�b�H4H���k��f)���E
��O�h0,�3䨵������g[�CdT�����wWW��8�66�l9����=5��q�$�Mv��~�Ȉ"'4cHcC�=�w���"��#���?ֲK��8,�3��D�¬�J��,)�6/0e�.`!E��A���β���3���ꎲ���o9�ZZDݦ�뚾b��i���8��0a�ž.w�Ʌv�r�09����lhcB��9�{���}�f�]%�Y��!��D�
[�t�Se�e��,��,#n�F�6⮯'`Ob�����1�ڎ�n��H�$�1�������cHN0%�RCNxκFNH��ekK%�R�	�JS�x~�H��r'~�A��Dz$��""Q�"(�������}nI��w�є�`�*�M�?�����@ax(s�1�&�8(+c{��:�rҸ���zN��{�a�w�>����rpW~F����4�{R3J���v6*Cf\l��@a�a�.q�����CE�| �X!CDB(H����|��ٿ�Ț) op����;�w���m5��{����8�z�W>��g��ঃ�C�,/�W����(\nXbeDv�\g0Y>��`���o����q2�w��� '}��Ȉ�#�<bDD8�N�" �1���G�=�gc���H����od�F��&�{�a+��ד#H�(�E�ۂ�ބ�m���\H$4�IԤ-�q�cn�ic��s;�La65���|���i{M'3�g*�	��&��V�XDYdD$�߄����vfΔ��m�ڍ��ի�]����v�̔���~�f?owA����q�D"B8�I��V"V3�ͣ�{#v�r����F�C��2��j���Q�lnLSM��=��_���#�J`n����b�8�������-��F��zg��p48}�8|�ܬ_1p����,�$c�'�f�/���YY����B1�7�&X^�W>D��;�;�n�Н���L��͈DH㈂�b�-�݇qC���v{BQ��!,>���q�)EvɊR���r:���	
Vm�2����b�Lu�� ��d����40�!��=D�yR��:�}�U9�Z�hDb*t����P\�&���iy9.�����)��c��)0M oi ���i�F!�~�>�����N��ߛߞΑ�=�":󠓪���١H� �a�%�^#��s���D��� h֙�!d�c�
1�6���u �ȋ��t<y
`�1����&�i"e;���G���ϯַk�����Y��A $��A!R*B���X�dePͣ��>��|q�.i�W���C��}�����?l{��qo��83gǍt�4VS�N���W�ǿWQȃgҬ�R�����<��C�-�%!���ͽ�5:��h��g��S}~ÿg�ũ:����ڽ���S,\�/�(�w{8g-�pFȲ`�Q�ްrS��_m�黨%|�qJ$d��=�Ua��f�O`&0�%���k-�s㚚���{��>�l�k�Y4Zk��|k����,p���?�7���ǆ~^<~������i�Fp�⊏~�N"����*?QmqU�vJ���ƌM��zz�g$Y�Y����Я�ϥKg��Y���&�z�Mt0{L��׆��Z��}��;��s���%٣������>)4�2���ɒ֙��u�]g[a�kX��ִ���+��\�j��e٧����V�Zִ:M��7NcUu�h�ڞj�]�Z��Zֵ�kwZֵ�bէ�m��.��Z�:��"(�L�ѭZS���+:�zW[<.�*�t��f�6�kj��u˕ڲ��b��I�Zֶ��ɓ?�����Rtff��L0f E�D0{3�i�5���i*��!ӥ�)	wF�FC�ы�H4r��цY"�N�%8�)N!��H�Ta���az7�8� ^MfZ�'�ƴ�lW�kQ�^�r�G7C<3��j4�t��'��w�<{�b���"�i��0��S��1���h���bB�
3�(��#��m 7��)�޶C��D7��֠��g�0ݦ��)��P����<�u����VVa� �Gp�\ֶl��tt�1x�l65��lg��pa�F�pV��T�A�����Ã�1�lv������B��ߜ�R�`Ϯо��\�Nlj�ta��ܐ�K,71/$7F�&�ԺED�Q�������@��i#b����y�`� i`r�����m]&S^"9!-��1���.�E^ən�����魋]#3�d�:��i�?~��M��yQR.�)�K5�vC߸�z;ֶ�B�ť�osER�B�I�I�t��BMԀ�k�ؚ��
�3�b���"hv�J���YM��ӿ}�D4��N ��������R�g�]���5����s��:���� @�Pd���@���	���.�p1c�;Ne�{���wr�F�"a1�#^��W�{����W�4Dq��s�/1�rA�c�\.1��b#Yoj;�n(�:����~�s?CĮ) �c]�9Ͳut�d�a3)H'�)�U���1����;9,k���YI���^B�Gt;�w��#E��~��B
�6}�������c1��%cL���W0�LB�`������u�s�&��M����tf<01��C��/��[�||F[F��E����B��9�N}��M�6���}r���3{���Mh�I$�K��u�8������6�
�h4�����"żv�y8r�F&v�*���||L	��Ze}B��E5���4��h��t~��"`4��y�O��f;rm����}��H	�����tT�"f �8'�4�#�{���@Ҧ���y;�1��68Q;�9��a�
�#��9�$XHFH��T}�,lac6:@������ey;Z$��P�����!�j&�ަ5:�Ǡ.��Z�k�����	_ْ�z�����(���^�$'��І�Yl�IfkHh�њ �_�Ҁ��m�� �=�X�"*F�
;���T��t�IJ��.�i�G~��,��#����Z޿	�{���{�#��Ŷ&@�L�1Q�	�[�ۆ*)�����x�)�^������\���RLLA��XǦR-J<�áDH��!pbo'l={��"/q�=�Fu�K$��b�g}	J�BbDp���!B�b3�c�݅�@̥M�5� �2�!
�%iZȱF��HO���D�j���0z����@�DՈ������"4pI����j���\��y(�Tl��w{����z(�X�R��q�`�)�te����*�ډ���k���kC�l��� ]�T!rĿbxcy��t1:C	(�JC�[G��w�C��ʉ>��n"Cт�@{�}�̡H���ㄮ��P��s�~|��C
��9���ښR�ΐ�M�o$1��GPB��N&��6;��<����� v�QkFM��bΔ,�X��}�
� �Fjc���=s������7߽>p#a��;�7#���-s�|�	��p�4�C�ג��j$=:����{��w�\�.0-4����]w�j�-&�6���s�Q�(�Ml�v����
R*�KY(�g,����@N9FZ�ے��O��������E�8c����GQ���*,��o��;��.O���Mof��M�d���$n�M��F�2+B"F��~��8��8����������Z9���b>��w�������k��dCٵ��{?�_�}�_V�[X;����!�(�x����
?[b(�ֳ���8�4�0�g�1���ߴrx݇a�x�=�W�o�)�j�f��wG!9
�)шl[���р�>TJf]Q�|��7Lyf����o~;w�c�����5�M��>���9�d7�<C���g��C�3��㦙���&��;2���~>u�?�_Y��#�L�I�զ{����D�q��(<Yԏ��~���Q�}����2A㒺�z6w��z��,*��.7��z֑6B���ѷ4oE�i ~5��߫�ppI�;��#�3񢇈r�k�SF�/���4�q�ދ�T(�!�|/ɒ��8E#x�c��8wC4kT��%�/~���>5����l�7���,p��72�-�º��I(� ����~,�d��T@�T������U�UU��.K��b,5�Ф
`�HcJS	
y"t"b8N�!yE�G�&Ɔ�
�t�ԂJj�Ϧ�Izݵ�۸��;;�%�t)nhA�4æ�k<.]f��v�G�n���ݹu�R���
� �Me� 3J��餘�gm��r�YTz�k����w/X��v�i�Z4Y���)L@�0R	�a:S� ���lt ���`�P��%4e��Zȑ.�K�t�E�Ϯks�����Z6�{�۳j���I�gL:���ZY*��kDi�F1K�gM٭��L��v1�v�v)�f{w+w8��"SLP�1�a��$1��9"[4e#���軍�$JA,J6$n,�!\%�P�x��HH��܋�ݚK�<�F1N7�>(�{�8H���h�ע�\7�Ʌ+��b��6��qZ�si��n^w;��D���)n[�)f��G
D��ʳnؕ��Ռa��C�Z��!�F�bq�{
%R�"c	�1�Q!�0Q;��?��C�>���Ƴ�����
t�#+?4iCF!i���1������~.��:.�l�����x�Xga��	�l� c�R���MA,�asM�З<f���<sb��3����cчHB���,z'31�,e���Z_e�����:Sz�]��M#P(�M]�3d9�t�J���6Q0��2������4C��	��6`��ц��D��5t��W�kX��1	b�ʪ��u�˲/w�G ��$!6p�����1��6�����ϩ/�ݶ��e�Cy(���'4%qyM�˦3N�ɬآ�s�,W]���c)��`��V�ܵ��t�Ś��3�R����)1,p�$tw2B&8S/z3>�a��BL���D�@Hy�F��ȝ&��T0I(���c(�tqs�\���+%��!9PР�1IiO<��0z���'1�NJ�GT���y�H����iU�s�,-"�:��|LL��#ݞ�ϲ��_1ozOOzȳ^I!��<B�GR�3��q����gC��9�'0�OZ�����<��������y3L$DD���� �4�Ǣ�X�~��T�֮���I�¦��\����7�����}0o;�����S5����td�҉�Bh��J$�nŦBS5�����8�����Tz��aLMD1�����d1���<A�A ���0�H��)	N2��L?\�v��F�1kE�9ޕ����Z���i�{�b���pw���>��G5�s�0�b��	9B��!I2Ld!L��e�[�>��oIE��c2���C�J��5]�|���
�/�>hA���$���\��v�On.Vմ�{Uu�]��ʸv�q�1����)Dy2Y���2RZ�Mi�c�Gw�oJ!����I<�c|?!��羲��q�!%P�D�妖��/�|�*���0���������6�4�5ʏ}�EZ�$mF蟽��������􄍿��Cج͟�H9��c��)�6��a1�!/t�yc�Z����)�]���;�'xYr��Ba8D��"��������p@��N���D
Q���>�8���!�	"]tD�^���v4zkH�R�H�&7C��Ŭ�!�f�<�'3�5(�$sAJHz�<ĉHR��$��B3&Cb&!L9Kh$y��:����2L[8�"Ի}�a��Ź��wS�@��ѵ�X��ϑ>av��}>0��M��#Z���g8b�vgR�^F��
S�5Q�`��i9���$
�5_�(�Χ�R��ҰD�BՅFZ~y��N��8��|�ĳ�q��e9QŤw�Ϥ�@�ڼ�G�栨0�}���k�d��U�680dm��7��iDi�ԓrN�q�n��ï�{_b8A�*���Dm�P����Q��J$+
��7p�]�u�V�	Џ������|�)�/��f& T|�D��ؼ�(����X��m���:7�����ïϟ=K��'����N�jꐦi���a���s۝�w���i�x��\�ޓ�DD�\C"��ih��-͇�8�	ߧ�?;sm��V���;�Siws�ݎ�ɶu���6:}�/�п��(���!'��x�ж	�B�
�d��[pt�
���~�р���&L+�d���o&kp����CQ iE�Z^z�,�2�6��l;�?��Gs�
{��O��h~���!͜�!Q��GΡ���>􅲿�� ���9�? _O�s.9�@��k��
�BB�`���e|�;��ݴ�G���#ۑ��0�:1�#��1Aj�u)��]R5FG���p����'�1����n�����M�^�p��ۚ����2�1�I""�����;����ЄCAH)"	�<z������D	 k�d�|0cʣ�=��f.cc�K�4!�~�!��A�N�D��&��:
��|Ld-0&�5�_86� !�a60�w��8�UG����~��e��kWt]�y�.����4����F�*�����i2��;�9�9��o��"9U<�H��(Ȣ�H#"B(	� (w(��nP0�?G��)�}x9���䄄`!�b�
�='��^^�@�aV��9�= RQc��Uu\>jb1o��?��W��?	wA�o�ӱy�BK�%c{!Q79��b�`�Kw�Lh#i�-J���H�Ѡ���}��\�������F5y�w������<�OS���:��4�܁�������֚lӌdf��O�+Dq����,@��Té��-�##�cDI �:���q�	ʆJ],�D�$#�A6-��j�4ș���:O�i��I�E�|H.L���0���ݞR�r�#���$2{齳h�:21�N�m�O��h�+���"P|!G��f˳�N�F#�2lh����g�)�߳3J���������<LKc��a��q�i��E����80Za��<����#G��h͌�6�;.�����Plh��=���11W��KF�ߍ%�y�������b�+ј}�9�h��>8���zsd8>l]u�/�cA�B���q��2���p�tz���>*c>x85�E��/	<��(�t�>��ִw㱞C4������c�,��+�Te��U��Ü.� �se���u�����D�p�£!>:VX���5�6�:Bҝݏ�Ґ��c�2聢ǹ��R�h�'w�g3zi�3����B�,��{n����_i���'�$B��QC&���)�; ��D]A:��m�h�f/p�r�d�<#�1q��K������ű�'�.�U����'����,!!B
��d��!!	\�Rp�v�{�ݶ�����c���kZֳ$N�5Tu�WY��ӳi�s�k[mkZֵ����kZ�v�V��e֮�j��Y�k�*�ֶu,�=��v���3S�nl��Cm��C1�I͔�Y9�Z��b�r�ЬBIB���_&���K�$я5��^.�)�C�4S\�M�q�;��k7���v[����X3k4R�I!��mr�k���k5|o����a�a�#�B��
��C���(_|��M"�w�{ń�C�$atO��=�X�h⾳2������D���b�5gs
ᔦ#k��9��L&�a��!���Ul�g�@UeS,,�~�B߽3�B&��e�;��!(|V	��Vs�EQe�=M-�����g�HDCD�.�r?�Ž�kgQĹ�F�hU!P6��$!!U��"
a:!Rr �c��Ix2�=Z)O��w߾��C�����3-�h�#4��FRr��(�ʐm�!
i-5Z����n��_2����lj���9��Z@��+�s�l���������;��O�Ư���ڻB��ٝu��3���Y��v�FbM��vIg��AE�J�~�u!2P� �	RDu�.�#
G����L��O|.[�6?p������I�9�LJHHR�SJ����oΩ��xO-��e7D����B.~��/O�~q"aM�n��_~�bh���n}c���A�\��q,��pVH�u�l��(��N68�q/;̝��*�5��m��3˵	�0�n�oa�ۧ�U�7+���v0����F��p��3��,%(�M�t�GG��GS"a1Ja���"��T���@T�C��Ȣ�w��<�8G���£�M9!�u#f�b		6&a�)J@hh����~�kȱ�D�/�|/�]��({���.sJ�}~��������Ik�C��#y�{�ʦ�h���1��İ�!y��f�9C8�Y�"(0�?5�&�1@B��220)88�~�T�I�7娜�(i�ZMA�"I����s��T3\oo���ѽm����F��y�?��������'�H�AVv��Hg\8$�䝰��!��v�u�r�;��V���x���Ɔ��䍉��M!*0c��D	6$��б�1k�߿j�29J4y�_/�CaF�9���%m��}˳K�㴙&���DI�CcrB4��uHS�����7�E{�j�4nm_�~����d�6�;�sM�x&"���|����gI��)�m<��ݝ��� ���)l��d�$T�;�|�� �AA�!���"������Xpk����8�.�ؿ�m+�?���[�FM�ba���d��i�c���q�	~�����D����>�k�A�Էy���D5Sp����шa����e����&�y	%��$�;
\&�z�& ��!����$�����g(�y��.�b#H�&56�Љ����m4Y��-���:��;�E�D�8�/!��S�؝;
C,$��$�L	�^%�1��Fǌ�9���I�!]NFr�2B|,���#�$ceN`�<0r��f�F�|�f{�0(�[U�_8P��q�P��_���h7@����l09Ν���f�u2�?8���-
j<1;�{���ݐ��bG	��A��15i���y�!t0#���Qh��E�hG~���45��������n���CP-)��a4����$��M��X%l��DPͣ�y��.��?8���ߞ�ڄ7R��D��d�h�)A�qFQs����9T�D46)c�(��|ޓF��@�B�`�H0�B0�ȩ2��!#:0��p��!"��WG��hh�@wP}H�/�<�á��m{�;	+�\n4%�P[��e�y'"0#|��ICi,5��C
	""���P����a�4�&�j�Q� rg�b%�a�CcI���m&�7���%yS�ֺ�Zƶ��\���v��J@�$`E+�6 �[��|#�B=x�%L�kc����s.�+�G�߼������{�,�&�'��9�vY�8�
T�5!1
YaJm �i��l6�	�^�o����#v����2"5�1."��}�� �ک{�O�D}Vc�X�rUJ���n&�����	����	�������?�>�c�1$��I$�I	 �H�

*%p�)��TOg��#@aB�"i UL!߰�K��CX�H9X�����%-�$HA�QqUPϳ
��D�����
���;X�X�b"�(��H�=�PP5EPS��&�� `I�⠢�d;�� (�����"�"��L�`Le�(��
��
ؐ� -�
����q-��2 G�H�q�(� �8`�",�0�:0�����LVEDB��M`��v8��Ł����t�}���W�0;��D�?�
(��TAD	BAQaTOA��>�C����U߫�;߷����=�ٕp�������_�5 ���ڇg�?�8����8�y��		<���g�Rz������O|�Z��p)����:�����^����z�KD�'�\<�����hJ~��'s	"WD�|���,ɑ����O���>xd�vz��@�h����Y�$�!��o�|G|��?���̟��E_CͿ?��PEQ+�"���_�~�~E8/�����~�����+�������Z�=h�k��s��T�������{��5!��?B��*|=����BЋ��?ϺEQ'�E>!g��H��\��������$��>��
�D�&��C�$�K/���V
pu�܂;І1��E�K�46�H�ظ����.��������S�y���X��!؇��>ߏ|>�O���t`�H����e eo-> ]�@�O��y��I��Q {�T�g׬i SΒ���F�ڔ$bF@/<*<<�r��"�
���"�� A��A�d� $FIDIHA�E	 �!1FaE�H@@$�YBB@IA���Ā���Ȃ�  �A���*���# �H� $�!*�*Ă!"�1H HH$�1 ńa,�aED�E�Q���A��YDE�dE�BE�dX�Y!!@A�I�P�@d�AW�{����xxD@�D	��@��$���X0$���2 
��p� p�r�"�� $��(BB�Y D$A�Q$Pb�A� "@YH1@��$D�$0@���REP�$H�RAUPbE�FdE�@$B ��bD�A� �$ � Ȳ# �S��P�x���Q"A��! 0`Ȅ��*��"�$� 1 H�#���`H$��A��H�`2���a1`ȱ H��H�H�#�H��A�� H�A�� H��`��H�H$��H ,���H*"(� ��* ,���"A�� H1"���H�@�RD�#E��	 ȩH D�$R! H�A��##0aHȰd,�����('<�"�B$V$"���	F"�'(����(''=ȣ A��� HA� DbE�9�{�ND�D�S�^�9^C��PND吃 �"E�B)@"@� $� B@ �d�Q @dP�d@b@�1E��XP���(��ā"A�H�  ��2*H #H�B �0"H(H+ � �ȧs��<�)Ȃ�	�$ h��a!@D��U@(H��[0
�&1�@
� �����"��$TN!}��!��bc= =�Q������h�I������~�O��
��h ����`�w�}�O��V���
=���tv�~H9E���#ϣ>"|�������~�� �c�>X!���?��]	�W��>����y�D�?L~���T�?�����!���}���h�*&	'�	N�����޽m4��}�}����;��D=��QЗ�����e����:��I�	�����i��G�� O�`��v�8��H�����:{�:�|
�,|@���>���q�����>����=Y���B(������tI	"�¿"�-������ٺ��Q>�^�o��oh���z!�_�A��I���>���z@U����ED��h�?�w�)��&Q��A �QhB��6r?Ǡ�t�hAC�nAOا��)AD�������1$ P�(Q�
�\>�_��&F��*�����O��-t.��҂�b���$L1��=��h ���yb���P��bA�0��}x�l��8���0A��'`��/A ���
!yC4�@aZ��2���Gb��qS�A�[EQ ��o�Ɣ�k������?!�ژ>��EQ=�~!�:?�ڿ�|�����g��� �������?�?��:��+׼~P>���@���}����B���U�"��?��¸{�>�>���{�_��]a$Q}��6N��bt��m��t.���c��p�"�c֧߂�}C=�	�W���"|&(�� D���#�����T_�0���*&w�$Mh����A݇�����@O�$�	���W�B�9N�=_F*�~>��}?w�菰��X�C�'��%}�}��֨�1�j��\����ȇ�:M���}��G��c�OP�E�~���J�R=�=t_����~��� {T�&m?��W��}A�"{QDTN/�:��r����:�,ZB��p�ZD�� ��A}4	���i��Y��I���!ߠ�.�	�����`�
��V7���cc��!`��b��(M���/����p'��T| �TOԬ4���Wᬣ�OX�R	��~���Bc��\_Z�J �'�Y�b} ���=�&��D?1��)H}��ä0���N�p�BӴ���'�??֟0�f>*1,dHX!�.0���"�d"l���?!�ȋ��rE8P�~�