BZh91AY&SYV�� �1߀Ryg����߰?���`N�r����l��E�OA��`@� ��A8�U	�p��ϣ)������f�f�C%��2[mkA��kIU`��F�v�0tN��4�v�c�����(l	`IA�[	��� RM:�R��S+�m���u�πM��SF� T 
@BUJ0 �   	��� �����&� � &   Jd4� 4� L�P��5PB�@h�2dh20&#L�	���� M&�C��h��h4�A "�I��0�##!�  4Y�6�1D�΂�zw������((�0A@ "(��A�<�<7�� N"#�Oh����Z��萙ť}�6v�j�щ��R�ҝMv,KP��^��J��-A��`��"_�EPJ�kS����,�%J�<�� "r��(g�~͈x���l��4D��3a'�f@�A+?+LK�����K�/�cӽ�l��
�^���e��ƀ��g����U���Qɩ���u</jG�e�&�43��:GB�ؐ�6���,ڕJ#ε�c��v�<	p������a n�>ؽ�"���Ӑ�*�lJ`�I�b�)Dm�W9��7b1��g��X܁%"��P-]3++���1�7�}T��@�c��6��F��������C�;���X����JE�3��8��v��k��6D�h��i�7Ll�Oy�yCs2'����V(3���W���P��b��g 9���/��((���{�!q��K=�^m�E�h��6�>��#�1:�y�>�ryX��D=H[x��j�:��:��}�C+E�h"C>�@Ԙkk�2mN���0���|�{8�xyy��%�)D�vr��ù�D�N���5A֫���i�j��r�^<|�����0Pa���@C~��z|9�vI�&����K�oO������x�"�5yy���	~�!!�����Y
4׋5��(V�o�����FuP��+*7Z�{�{5�i��K�yNcB��Y�d��RyψHJ϶���\@" Q�	%-�;���	K³�c�N���U��x`B,�aX|T��0�	xE4�z��)�y�rՖ��xfb`� lBȦ��C/�\�R��8���Cmm�C�>�t7PJ�o������AY��1�O����䑪�rS�.��h�@]�+� $"�2�2X���h���1 ��Q���F 9�
����G5�Mx$>�Jr=�%��'�/3q ���V}�����9���w̭��2�!B"��`fPM�wg�2 �J�:�E�!
�����K�3@�$���v�;A�U�����Ro4$�5�	�M۠+�/�%�q �X�EV
��Rݵ��q�t�;K��
n�W6�H����!U�^�E��`�WA�W9��x![T4��5p�)�/#��i���'Z��Bڷ�K�Eou@�ᘶnc����\db�2���	���+6����,�E�"ƃ��qvPT�z;�!*��䟛Z���o��͞�H��*�l
����Ko��\�龜l��͠��M���di.7�/(;n�/���^=��[�y��<<��y�/��M�������y�9�9�+�9�g,��zm<�&t|����=���/v���<}3���_E�9�5��λ�q�$��Mo9��'<烞s�w�7����:g<�3�s�o:g=絧9�<�Y�9�g9�<磞s���7^�u=ٜ���Y�M�{�wwo9$�Ι����\�N��y�s���<\�s�/:��s�9��ٯu���s��C����˂&&Cp$ �������v )S�_�3��.�N���Wa�JN����e��o)=ݘ�WIywwi^���{�w]<��m.��㧲%����R9�9�?�u[��m�W��a�3j�S_m2����0��3>;��:�s��>%룫w$�=�f�O��Τ���Ώ:�>�Zw�թ���V]��������7����߸ȟbt]?�m�I$%��.���ty\lp��A����͓:�mZ����Ӥ���d��}��VeJ�פ������y�9�n�s׃��wR������ˑ���׽p��ŖV�`ɏ{�|��o�=��d��I��$�M�/
�Ʀ]����QWgU͏^sΒI>��N#�j�$��C�vUt�8Vʩ4F�:���KT����vi�����p�nhg�H�[X��Z:�~Tr���rי:��Je�y�;s:�NvY��H�z��j��w]{%����;��p��E�k��=qR7>��*�HQo{o��7y�T1�CA;q�I�V�4�=$��(��̪��|�ט���	#Ǚ���y�i��ogwV(b��q���5������y�Y�|�e%�ŻΆ�T��ީz�u�˨�:�['<�Բ�`Zx���;5���0XE�)UҞ��V��g+�N� e�j�N�Y��i[y�n�ܭ]���$��]�y�܎r��wo���Of�ܒHdJ�`�O1��rH�v�(V�N�iP#s5��T4[je������篞��9�<��Z���M����l�n�g2��{��x��y�9�<��IΛ�q��u˭�{�M��zglV�7w71���s��{���X�7I�)�T�H�|}�{�ζۼOga����MYD�E"�M��j�hv_v>ל�{���u���v�^s�y�9�s�S���]�h{�f�)�����{:�{ikd�e5N�y�&I#��B��[��k��m�I�hma�[�t��Io5%� �1ͺ�Xa���j�9�r������w']��޼��I�T�����e&7"�G���aU�[�`}K�0��Ț��_�����"�8t0�h���~��˿�p��ǲ��]�
V���^�m�� �C[M�B�F̱�5݄?1���Ψ<���[����66p� �x<=��"@���Q�0��kٻ�
H$b �:ܹ��)�ҫ�����@DwXR�`(eV��r�t�G&���g^N�̲H! @���^0�����$�*l�ױ  �c��6�|7�Um���]t�&*�����%�=��:g����V/x�G��u�T�9�ͺ�[i��� :��j�M�COsT��
�\q,݉B�)c�	�� �!Rma'_&\:wJH�D��U���:��2��Vk���X[Vf;�կ� ?:�TH���ݽe� ��&5M4�q���>��G�X�����p�
� G��\�` IJ� p���w"��ܨ���S�G+�� ���os�ۣ�.U����=]�5�1{%�u g��Ӎ@�o�fpU��ۖ���JW���w>yi����;^
�T�wW@��2n����\�F&4L���E��R��O���%EA"�bD�3������
%gS �$]��<�6mr�'w�N�|�u���GZ��%�[nxź�&��]�%Ipͱ���p4���K�uƚ��d�[�� �`-8�k+4R�#
�֓*f���ƛ6e�s��Xl�͖]	��hw&��rϰ��s�'�=;�~G��̺)�Cc� ��:�b" �S�m��B-Dͩ
n�D��L��$~͙ ��d��s�V��M�.�'�$5_� 5�{�FhdqAJ����L�B�1bc��h�H�k�CW���|��C`H�g��+1.��8�
�Z�cI�VY�>mί|>��M;�����iv$lo�M$��R�Ŋ`9��3{�&��D��H.��)s���{ީ\��k�GZt���j0��~?��|s�T���AD�h�\�x���lR.�v8��?(���=���<<�b�������[ʜ[
h��e�Q�$P�9<x��z�ىfߘq�lE�v���T��,5,���t�@
����)��	��X�Q���y3��fި:ub{�D��JJ3��˦rY�\���U���a<�<��K��e�3Q�4�ě�MMds���.���;��7�i�xU��8��O98�&�����Y|���n)a�V�q�#7P�h\��$�e�o
�#�^��'T�F��t���i�r�Ӵ�o,ۜ����B��;��e[�����_m[^A	�l}XAXٝ`)��
͜�[�bV8�v� �@Vi�)!�b�E�/JEU��4�pJ��nx�.2��K�0��K;�m�"]}d
���՜��b�/�b�c��$����;��1���О���*�d���&��T������晙�kZ�-mYZխم�hk���Ɍ�CdC*�WR�Q�4�u���Ҵֺ��f��f �k͛����6���6<�ܚ�H �o����_9 Z�s�21�$�R���5����661c��QC3EB�5$��n���b\9�eﺮ���T[�t��,L�jr��{T& o���S,s@׸�pH�$�$'VI��|����n&��i��ͪ�*�ONrI�8�UTe�/4���|�+Ҧ�7��%����$�m��C�gZ�Je�R��LG]��l����B�o]0�^�8 7D�A���sȨtl!�o�l����ջ�j�ؾZn]TeUII$DX�2ɦ�f����[��E�����Js�Q�-�3�[��!��s�����S��͝��;���Ls��}���pv�u�X)�w�.�BA�����$��9;�tC$�T����j>�מo��d�j3꣙�h�G��*��,F�K���.�{����4FD$aF�DY#R��B#�Q0Rf4E�yG�R"�x���KVg�kH۱��Q��V�����̔�2��؄��9���������g�,EƗj��*ۣ֔�xNs�䤀B�YR���p�CP�/�[@�%x,��J)�:�Ap{Hf8��t��F��FO��E h`FdC�>��I�tH�s��g~m����]�i�噮5�m6.�J��a�� !�ЭMT�h�E� �9m#L�rov��V꽲���1�hMn��Q����I�h
@ v|��G:wͻ��-��� Cδ�I"uL|�sv� f�����LD�..�����-�� �_�Nƣ�l�m��b�|]�s�ߔB)���+�%6��7���C�3�/���`dE���vVP�{1���F����D�)�������+~�����\�y	�o��uJ��DV�ɕ�^�`����zy�g'���ܗ�L�߇�4f7Hb:"�>�J3:@�Gx�s�#{���3��w��{���Vyܔ�'�<��j����suW)M��JF�o�q@X���qd�-@�J��fV�n���u�V�{�%8O8u�����0�6����j��"����9�i��B�i�^3-0�)h�BP��YcC����s�)z3��E3n�	�&K(]�[V�]��ku]�%mj͛r�.,���Ũ���g|���8�������@ �}B����%U�҄�uZ��bhNzFގrs���#�{1{�qm�y�����M�ړm.��W��Փۣn��EY�Y�cp{�����3�K����fb\u�B�8����-a(��Gh�WCv�Vp�"��� .�9E��'�j6��@,�%T]�C�pf�1n%�p3�Y¤��W���tPYa�s!�G�ҙ���<(R"�5���h��i�@:��e��'Ͽ	}3&9�	�^�f�L-D�u��Q��K�j袃1s �<�P
)捈�tW��]BQ�Z��e�t���`u��ӟ}$h0G��ͧ���0�ǀX0\DX���¨���޷w�j��(��B��D�0�x�tG��m]g�(�0��%�A���k��@�y|E@hPqA#�ڎ.Ԙ��:�(G}��Ǔ�7�>(|ӂԕH%j�@�OOv��|�\=��"������l*�{k�2-�	��VdwǶn�9�F������w�Oz*u�j��B��`�dUgֻ�{s� ��	����9χ9$�Y#��ɭ�$<}tM���v,�2�v����Hެ�{��B�=j�xzl�NCu�-�ǒ�d��6ػ;`�G�
	$�2��bqZ��!��3�C���Gq)!�6�=ǳs���nZp�p�hK,=&�I��be�Pj�7Ƒ� #7l]��L)I��"#uɡ�Ѫ,�kE���a���q�����E'�!�h=."&cz=8'g;��82�f�(�ag��6_U�|�Hh<�8��.���N�h�Kd4��	F��Q�*���w
��}�1�
 #@b8��5m9�Qh�@� �4��K\�{$s��+����9�H�Gs#���fy}�v��F�;����f��ºN�QE���M���|��~�e~n宛mW]�kW���n�jմi�7mR&�B"m%��c�2@R���u�b�`m4��Q�W��K]�����U����s������$T��s�pȧ����qp�_M�P0(�� {+�TG��f���A.y�M�Z��"
gL�`�៹խ���Ȭqk)�ɂ1�$ P1���"* f�R��:$�M�w"���k?cq���u�:kcQ�'��J1귍u<��l�"汙�%ق�����s�<�`�nj��x3Q�"��MFu>�Ab�0)̋��R|����hO�G�Ջtxɦ�\�2Pʁ'�Ȑ�$����}�uF�a�@Tҁ��3LA\�Y�M���"ǰ�"��`9��$<�Bw��gN@�����I}\��d��Uw�f� ��֘z_F`BD@'Y�Dr:�ꨁ��{��2::��޷�=!�����ho���1v2�⧇���*K��ywbǶ��Up���u�䛚�_��s�������Z�uv���*����ٙ'���_�y�}�����+<[r�a���=��0�@L��ř�¾�"�?��T����Kt�����<���G�ҴMV�"Ca�K4��Ά�����~���u�J�7E��U{̀`\&n�վg�r������T3D���=`�h�{Tb����G���3Ζ|��W,��ԓv�"sY����= _%X�ť"�J3C"}�4��L�7a�Gs�����BD��*�.����'����O�X��P�]�.�a�3�}&����(�!q�A�sug{ȼv DDD��M�N�a j���R�v�S�>�A&N��	JU6���k���lT���@�%����E��@O�¡���'P"�R�=
&�7A:&�9��4�"�r�@8�	 �]�n�<��� �e�.�f�9]I�7p��\骪JX��pvu�k[dRGT���xn��uu���嵗6f�ݲ���!x唤ٺk�`�ѻ�W:��-�یLV;k-HX��m�\��<�YO`�|o�b!�7�� ��ŗYP�Nu���!j�T��� �Î�z�����9�I�sxzm�8�h�fAYe�*j)vtۖ0�ŝ��=>�A�	!��ȤsЄ��s��m��a���P	�o�9>�=o�f�p]�g����@5�� P �J���ÈTA���\	�����a��*������*<�vT0U��x0`�P�2}�`��i�؊wB��|g��51,׵	��uF���ξ�����)��WZ�cƃ�U�=6���t(kݵcX$J1s���b��B@��eU{<Ě��O�9p�1��$��/')ȿ���Y��3� �V
ᤩ�N1��Ō�o�s�s�-#A+>�\���݀#>�2q;�Y�ҙ߸��b����|�@Ոg�A!a�zg�ڃ�k�Hw�A���&�	V��z�1�#��#��\�ߌ�޶��oEWRa�o��B���"���U�w�p��)]h7D0��\��x
B�K���a<�7�~�N腪�A����T��t�g�΄�i��+}��uy�_�������0-+c%�mf�	�������u4�X�O�2����$�>�ϡ�ք���Td$i7��}�];�:9j
�\� �(��xgu'�C@���%(k ����P�ǖRЎ�t ��- N�X�4e�Q�L�̶��s���eu�(�n-V��딻���ą���D��n��Ɋ�*�hn&.�<��ʐz�vg��S��2�]��b �b���:^[�#�&"!�K���\ֶ�M�[�[]�����Wf4L�efv���d�H8�th8�L�:Q`k�^ ����V�Bݝ�����Eel�^S��N�R����;�LE"�!I <ח��իX��Z�Tȑ$����$ �q _=�gןv�y9�~��{��ͱ�U�4�EA��%+�7=�@�W�w��Ϸ��:�up��7ۙL�Q(L�g���
�N=CЅ��.�y�� ���ӈ0S���D�b]��{?wm��X�\XjY��f��Yn�/������T>�{�/Ϻk������A	�wc���H"q��$�α,��
83��H sˍ�GY�H��,�c�X�w�+OFB�`�@O���]�o��LD`x�HPRb��1��5F����90 %��nM*B�`inؚ5���<��{�+P�d˒�(��
��B�#9 8@���jH4��29��%���{�����os����a����4�KM�q.C @�<�EZN��5�W|Y��8Ȅe{ب�f���5��b"��Q%�%����;����≀nsܩ7�G}������f�+��O�
���3����%z��]nY�o��(���'52(��@U{�ʒ �ϗ�o�-"��������Mu�+YJ��"�ىo����m��ϛ~�<�ʱf�rd��Be_�B2�jG��xV���{ؿB�m��'Ԟ�#��v��������œ.���՝�3&�!��I���S��wσV�vr�
Q[l��F��^h�naҘu�Q�x�Kmˉ���,٬��S)��F ��͡��LG�h)V�d���\ifۖ�1P̚��#��D4cf�?���4?M����[[�ʦ.��n��xy�+R�n�����Ω�d�`_P�u��&�C�X7J��u׊�X!����4DW��Z\�ӕB�7�E*�ϻ�l�ɜˢ���@��J��"�eOF���$y���X�Ƞ�=СNЉ�+�������N>���L�F!VΘ��U�b�M���(Kq� %w�fM����XO	�ν���$��W����MVU�WQSY�$��ws�Ͽm��zP�B�HBMړ����7�B��O:����\�WEB�s��}p��s.%YxUp�IY����X!��W��Ws�Q�	��,Us��;�0¤�"�=�W��>��R�#ěb ���y�o�d&p,�o��6���!`(7x9�P��á�7D�H�|� ��\�Ş	N��A�]��ψYY�Ds;��:�y�߹�_������Q���&aD!�;���6�z���Ó1�o`�#"�&M;�e5�r9f��f���O�����(�3lJdl����4��^*�`��_�+�z���:H��S0n�HUA��=�A����!Ҁ�D
��@1]�8]�<�@�nsMfL��q
;�0��f#���� ���TK�����)j}s>t`W���i
	����-�f��7�9��l�<0F����^w���,Wr��y�h0��rsî�'�������mm���v�k[�Wj֭[a�XF��H2���0XR�J�5r��B!��2U�3jm�p�:��t�.3jխ�V
ʹN�"6u\�ޚ�*�6�5���	�ҍdvH����A&��f�"\��7-�Q��_(��P�"{x��{q�a!M�0Y���'{�&tlQ=���!��X�9��je`�\	;�t�z ��I*�_a�H^"_}�$�^��o�ȅ��9�>4�9�E�G��A��Y����K��ɂ�0��Y�Vw�Np:��^����!��#�nvj/�eyܩ�ho��ub,ȁ ��	�q��6n
CYi��g�54s�f������*t0���V*1� �:dI���9Sy��x���2.�=(Pkz�BDՏB�P�3`�"�n�3�4k(8���Uj��l�[��������x�b�H�]�H$!��;}K��Q��6 U�p��C�c�ɐ;�Bu_O"ի�n����f�Z�x�`)�9t�4����^|�3,�Ci`_��w??:��|H@��15W�A�yq��w*ñsB!��;����ۈvH��	�2����I�;ą�R�I�A'K�x�AF	�����Bo�WG�*<U3

  R��}��v7��/u����E!w�ޗ2�u�d�H�9�bC�>�;�]s";
B
DԼv��7K��	rlO}��y����*��@�u��-[��3�sd�5y�p�9��")s�1pO #PH��S+ˋ���*���:Ρ�� ��K٣��Y�Q��<��;hH��M@K.��  T>��uW5�e�O%B��zns�Ɏs��|)߿����hWd������&�p ��Sٺ�J���mf�dm�v�t�6���s\Mu��u� &#\F�&m��f�aM�Ԅm�.�V���b1`��˴�M[o�?'s�r�i�.l=P���[`m��2I!5��{��WGd�����b�%�F^J�j���ee�Nv��f������h�����H�(&�p��sp����ATQ�7�b��-��BIh��1L�6�T�b��5y��A��*q�d�c|X�����Hyz�~� B������Mg���#��-Ŵ��B�_8�r�A�"��)��� �j���ۯi.��?V����r�6�.P|�$g��lG{㡥$Z�vɢ��Kk&xS� L����wP�B��9�V���I����v"�ʖ�B�1H�:@�iw�f�2A��H|��2�n9孧պ�x��"Zo����w7� �����?<F���_�aC��fB�T���WQ��C#�U�����.z�H��[�f<4���^�{�*����r��}�����Ø35���k	�^[N�߽uy�_��3�A�5^�=Fi�� �_�p�왮`O�
:�^   ��ޢ@�ڇ"�fV��Y�5c�.�ɂX�<K�uҚ��0��	cr$O��ɾp���@�2>F�'7Ԇ�����z�gs��%�Y��	r��P���`������L�?7�{�@��4�m���"�$�+iż��R$L�Mlp�O��|��v+%��Xwġ�G�����蜓�u������mn��s[�km!��+�]J��V�Z�T��q���M�\�p�-0���e�ٹ1W[]�p�����غ��� U���PkF�V�[�@�r� ̗��&��@ +O7·�Z��.�px{�D|��6�����,ewtl52���hCF�y��\%�5�N��Q�j7��V���۬���O����>���/�zсm`m� �Y�\��T�ؾ�����}$��Ʈ�ml�+��J:.�!���m�4�Y�l�n��H_X�:n�U{�gRpױ��qT;ĩ�&2� ����ѽ�Ξ\l���<�	k<�x��ˏKI1P�4w;�*k���p�@�^ e� �ڡ=X�>���Ԓw���0� ".�?u�2�Z̿dGy=�o�����]Z��6Nl�KUk���Gr2!�]�b�@
M�l��z��_��TX�H�wx��W{/y����i��R,+&��K*[f�H���%�wY6�Ǿ����UVGQ�e�Ω�^��H�,��r$��z��;h_{���{����o��	����7;�Hъ5�6<������{��44���|p�J���
�P�{�7xf$�g����k}��#�U&%�b-m���۲5���u��ν�6X��T঑XF^GX�A1.�M=�D��Y���'�ffY\��Ėo�p�1�|�C��2RI!$�H��"�	R4|��EPM_r�5 ���
�Bÿ�g����à��h55����
Ȋ4D\D@����W�@C�J�D 7  �P��%�A0bR*�[��^<p��ApA�d;҃Ȳ ��v�肂� 
���E  ���@ 5
 ".,�a��,rr�6��E����Pv�T|�\$�x� `�MM�JH~��-=8l������p��?�ʊd��AFCɀ��Nc���(�J�1�A�?�V���gJwl?�An`�W�
�n�3���ӓ���I��&��j�=Lm�%N��h�[�?O�J�)x҆}Ζ�<偧� _�֢�%c@T��7%��p�8
(Jz��@"N������ �]a
$�`2Q]ń�v{�B��u��n�>A��"��Z<W�)e:����v��hە��q���X��3���P��x�EPI�!�I�ڶ��;`��Ȑ
���������yF<M�C�9�ew";Е[)XЖ�ռ[������ѣ�\�776nɄ���Y��pW���������5�I����٭)q�<���~����4���l�C��Ԁ�21E�Q� H9�8@� �B Ca�ElUV�H2(H����"�"����+"@� I	#	M�@�YE�DA $XEd$Q$Hő�$$cE��@��$D�d	�aA���2B$d$�!A#DId� ��c$r�Ð8 �!�� � a$�@���9�
� �� ���H�b�BD$dh*�H�$"�$�$��BH@$	���$$a	B0jH�H�H�FA�Xd"�I� ��#"��B�I B$@B  B!p$p' 2"H� �$��!���1�BB��Ȭ��! H1�$�H�@���!�#	B(H�����)B���BQ���/?W�� P�.x�#z�^� ���J(])��uCY�A�r��s����\Lފ�-�ѹ��8�io�y��� ͓��i�~�3�xt_�`ʻ{�������3~GkP��,"�%
��pj�z
�t�	x7�j]�
v/�\s�g�����jC�|��nK�F��ĽKí%��I/z���)��U�G'/Pb9�C�W� ���s���!	N������Ս�!�\:whz+5v����A5qb8�R	(<S�ܽ�J�܌+y�r9l��MX���.�֌11�X=B%����%���EPI��6�b�.����G��J�`3� ���q
��0��1�_5�@/yE�9B��R�B$҅H�*5v��<�p�VpD�q��,��z*����!MW���T8MА���p�)#"F(�K��(Q���E���dd���K!�� Zuim����F����R��6T5�D;������<s*K��� ��:�U֞A��߱��6��?,���{h2XsWiatr���#���<�*>�|�3��HzY0�nD��{��E�s�����������Ai�,LŮ��1<��b��ȳO�AA)�<lױ�`!�!R��B?�U�V��y�i��aA(����z��#}�߯*i����gQ������N�(S�Xj���m���"ҁ�O_"��<-v��m��}q�nb�NǊq�`�й14���~�qCH4L�	����V�W�5T���`̘=E����Mٷ��M�*�b�к5,�v�)H�UĮŢ�HUE�@��F������sAV���;ԙ�;֍d"V�a���M]��xYmMo�T0�p���6P��'ԱB㇘\�����P�������)�_\�#��M�>��q2���oa��>�Ka�]�;#��M4v'{3B�F��=C���S}JN�B$0zQ_�$����O����rE8P�V��